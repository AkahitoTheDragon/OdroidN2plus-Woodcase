            (     (                                  ������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         ���������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������   ���������������������������                                                                                       ������������������������������������������������������������������������                                                                              ���������������������������������������������������������������������������������������������������������������������������������������������������                                                                           ������������������������������������������������������������������������                                                                                          ���������������������������   ���������������������������������������������������������������������������������������   ���������������������������   ���������������������������������������������������������������������������������   ������������������������������������������������������������������������   ������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������   ������������������������������������������������������������������������   ������������������������������������������������������������������������������������   ���������������������������   ���������������������������������������������������������������������������������������   ���������������������������   ���������������������������������������������������������������������������������   ������������������������������������������������������������������������   ������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������   ������������������������������������������������������������������������   ������������������������������������������������������������������������������������   ���������������������������   ���������������������������������������������������������������������������������������   ���������������������������   ���������������������������������������������������������������������������������   ������������������������������������������������������������������������   ������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������   ������������������������������������������������������������������������   ������������������������������������������������������������������������������������   ���������������������������   ���������������������������������������������������������������                           ���������������������������                                                                                       ������������������������������������������������������������������������                                                                              ���������������������������������������������������������������������������������������������������������������������������������������������������                                                                           ������������������������������������������������������������������������                                                                                          ���������������������������                        ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ���������������������������������������������������������������������������������������������               ���������������������������                  ���������������������������                  ���������������������������                  ���������������������������                  ���������������������������                  ���������������������������               ������������������������������               ������������������������������               ������������������������������               ������������������������������               ���������������������������                  ���������������������������                  ���������������������������������������������������������������������������   ������������������������������������������   ���������������������������������������������������������������������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ������������������������������������������������������������������������������   ������������������������������������������                           ������������������������������������������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������������������������������������                        ������������������������������������������������������������������   ���������������������������������������������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������������������������������������   ���������������������������������������������������������������������������������������   ���������������������������������������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ������������������������������������������������������������   ���������������������������������������������������������������������������������������   ���������������������������������������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ������������������������������������������������������������   ���������������������������������������������������������������������������������������   ������������������������������������������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ������������������������������������������������������������   ���������������������������������������������������������������������������������������   ������������������������������������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������������������������������������������   ���������������������������������������������������������������                           ���������������������������������������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������������������������������������������                        ������������������������������������������   ���������������������������������������������������������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������������������������������������������������������������������   ������������������������������������������   ���������������������������������������������������������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ������������������������������������������������������������������������������������������   ������������������������������������������   ���������������������������������������������������������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ������������������������������������������������������������������������������������������   ������������������������������������������   ���������������������������������������������������������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ������������������������������������������������������������������������������������������   ������������������������������������������                           ���������������������������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ������������������������������������������������������������������������                        ������������������������������������������������������������������   ������������������������������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ������������������������������������������������������������������������   ���������������������������������������������������������������������������������������   ������������������������������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ������������������������������������������������������������������������   ���������������������������������������������������������������������������������������   ���������������������������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������������������������������������������������������   ���������������������������������������������������������������������������������������   ���������������������������������������������                  ���������������������������                  ���������������������������                  ���������������������������               ������������������������������               ������������������������������               ������������������������������               ���������������������������                  ���������������������������                  ���������������������������                  ���������������������������                  ���������������������������                  ���������������������������                  ���������������������������������������������������������������������������   ���������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������                           ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                        ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ���������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         ������������������   ������������������������������������������   ���������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������   ������������������������������������������   ���������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������   ������������������������������������������   ���������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         ������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ���������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         ������������������   ������������������������������������������   ���������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������   ������������������������������������������   ���������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         ������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         ���������������������   ������������������������������������������   ������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������   ������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������   ������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         ���������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         ���������������������   ������������������������������������������   ������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������   ������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������   ������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         ���������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������                        ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                           ���������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������   ������������������������������������������������               ���������������������������                  ���������������������������                  ���������������������������                  ���������������������������                  ���������������������������                  ���������������������������               ������������������������������               ������������������������������               ������������������������������               ���������������������������                  ���������������������������                  ���������������������������                  ���������������������������������������������������������������������������   ���������������������������������������������������������������������������������������   ������������������������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������������������������������������������������������   ���������������������������������������������������������������������������������������   ���������������������������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ������������������������������������������������������������������������   ���������������������������������������������������������������������������������������   ���������������������������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ������������������������������������������������������������������������   ������������������������������������������������������������������                        ���������������������������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������������������������������������������������                           ������������������������������������������   ���������������������������������������������������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������������������������������������������������������������������������   ������������������������������������������   ���������������������������������������������������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������������������������������������������������������������������   ������������������������������������������   ���������������������������������������������������������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������������������������������������������������������������������   ������������������������������������������                        ������������������������������������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������������������������������������������                           ���������������������������������������������������������������   ������������������������������������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������������������������������������������   ���������������������������������������������������������������������������������������   ���������������������������������������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ������������������������������������������������������������   ���������������������������������������������������������������������������������������   ���������������������������������������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������������������������������������   ���������������������������������������������������������������������������������������   ������������������������������������������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������������������������������������   ���������������������������������������������������������������������������������������   ������������������������������������������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������������������������������������   ������������������������������������������������������������������                        ������������������������������������������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������������������������������������                           ������������������������������������������   ������������������������������������������������������������������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������               ������������������������������               ������������������������������               ������������������������������               ���������������������������                  ���������������������������                  ���������������������������                  ���������������������������                  ���������������������������                  ���������������������������               ������������������������������               ������������������������������               ������������������������������               ������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������                        ���������������������������                                                                                       ���������������������������������������������������������������������������                                                                           ���������������������������������������������������������������������������������������������������������������������������������������������������                                                                              ������������������������������������������������������������������������                                                                                       ���������������������������                           ���������������������������������������������������������������   ���������������������������   ���������������������������������������������������������������������������������   ���������������������������������������������������������������������������   ���������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������   ������������������������������������������������������������������������   ���������������������������������������������������������������������������������   ���������������������������   ���������������������������������������������������������������������������������������   ���������������������������   ���������������������������������������������������������������������������������   ���������������������������������������������������������������������������   ���������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������   ������������������������������������������������������������������������   ���������������������������������������������������������������������������������   ���������������������������   ���������������������������������������������������������������������������������������   ���������������������������   ���������������������������������������������������������������������������������   ���������������������������������������������������������������������������   ���������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������   ������������������������������������������������������������������������   ���������������������������������������������������������������������������������   ���������������������������   ���������������������������������������������������������������������������������������   ���������������������������                                                                                       ���������������������������������������������������������������������������                                                                           ���������������������������������������������������������������������������������������������������������������������������������������������������                                                                              ������������������������������������������������������������������������                                                                                       ���������������������������   ���������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             ���������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������������������������������������������������   ������      ���������   ������   ���         ���   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������������������������������������������         ���      ������������   ������   ���   ���   ���   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������������������������������������������         ���      ���   ���������      ������   ���   ���      ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���      ���            ���������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������������������������������������������      ���      ������   ���������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������         ���   ������   ���������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ���������   ������   ���������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������������������������������������������                                                               ������������������������������                                                                                                                                                      ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������         ���         ������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������������������������������������������   ���������������������������������������������������������   ������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������������������������������������������   ���������������������������������������������������������   ������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                      ������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������������������������������������������   ���������������������������������������������������������   ������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������������   ������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������������������������������������������   ���������������������������������������������������������   ������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������������   ������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������������������������������������������   ���������������������������������������������������������   ������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������������   ������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������������������������������������������   ���������������������������������������������������������   ������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������������   ������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������������������������������������������   ���������������������������������������������������������   ������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������������   ������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������������������������������������������   ���������������������������������������������������������   ������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������      ������������������������������������������������   ������������������������������������������������������������������������������������������������   ������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������������������������������������������   ���������������������������������������������������������   ������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������      ������      ������������������������������������������   ������������������������������������������������������������������������������������������������   ������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������������������������������������������   ���������������������������������������������������������   ������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������      ������������������      ������������������������������������   ������������������������������������������������������������������������������������������������   ������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������������������������������������������   ���������������������������������������������������������   ������������������������������                                                                                                                                                      ���������������������������������������������������������������������������������������������������������������������������������������������      ������������������������������      ������������������������������   ������������������������������������������������������������������������������������������������   ������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������������������������������������������   ���������������������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ���������������������������   ������������������������������������������������������������������������������������������������   ������������������������������������������������������������������   ���������������������������                           ���������������������������������������������������������������������������������������                                                               ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������������   ������������������������   ������������������������������������������������������������������������������������������������   ������������������������������������������������������������������                           ���   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ������������������������   ������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������   ���   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������   ���   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������   ���   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������   ���   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������������������   ���������������������                                                                                                      ������������������������������������������������������������������������������������������   ���   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���                           ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                           ���������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������                     ������������������������               ������            ���������            ������������������������                        ���������������            ���������������               ���            ���������������������������������            ������������������            ������������                                       ���������������������������������������������������������������������������������   ���������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ������������������������������������                                    ���������������                                    ���������            ���������������������                              ������������            ������������                                 ���������������������������������            ���������������               ������������                                       ���������������������������         ������������������������������������������������   ���������������������������������   ���������������������������������������������������������������������                        ���������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ������������������������������������                                       ������������                                    ���������            ���������������������                                 ���������            ������������                                 ���������������������������������            ���������������               ������������                                       ���������������������������         ���������������������������������������������������            ���������            ���������������������������������������������������������������������                                 ���������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������               ������������                  ������               ������������            ���������            ������������������            ������������            ���������            ���������            ������������            ���������������������������������            ������������                  ���������������               ������������������������������������������������         ���������������������������������������������������������������         ���������������������������������������������������������������������������                                          ������������������������������������������������������������������������������������������������   ���������������������������                           ������������������������������               ������������������               ������            ���������������            ���������            ������������������            ���������������            ������            ���������            ������������            ���������������������������������            ������������                  ���������������������               ������������������������������������������         ������������������������������������������������������������������������������������������������������������������������������������������������            ������������������������            ���������������������������������������������������������������������������������������������                           ���   ������������������������������������������������������               ���������������������               ���            ���������������            ���������            ���������������               ���������������            ������            ������               ������������            ���������������������������������            ���������                     ������������������������               ���������������������������������������         ���������������������������������������������������������������������������������������������������������������������������������������������         ���������������������������������            ������������������������������������������������������������������������������������������������������������������   ���   ������������������������������������������������������            ������������������������               ���            ���������������            ���������            ������������������            ���������������            ������            ������               ������������            ���������������������������������            ���������                     ���������������������������               ������������������                                             ������������������������������������������������������������������������������������������������������������������������            ������������������������������������         ������������������������������������������������������������������������������������������������������������������   ���   ������������������������������������������������������            ������������������������               ���            ���������������            ���������            ������������������            ������������               ������            ������               ������������            ���������������������������������            ������                        ������������������������������               ���������������                                             ������������������������������������������������������������������������������������������������������������������������         ���������������������������������������            ���������������������������������������������������������������������������������������������������������������   ���   ������������������������������������������������������            ������������������������               ���               ������������            ���������               ���������������            ������������            ���������            ���������            ������������            ���������������������������������            ������         ���            ���������������������������������            ���������������                                             ������������������������������������������������������������������������������������������������������������������������         ������������������������������������������         ���������������������������������������������������������������������������������������������������������������   ���   ������������������������������������������������������               ���������������������               ������                  ���               ���������                           ������            ������               ���������            ���������                  ���               ���������������������������������            ���            ���            ���������������������������������               ������������������������������         ������������������������������������������������������������������������������������������������������������������������������������������      ���������������������      ������������������         ���������������������������������������������������������������������������������������������������������������   ���   ������������������������������������������������������               ������������������               ������������                                 ���������                           ������                              ������������            ������������                                 ���������������������������������                        ������            ������������������������������������            ������������������������������         ������������������������������������������������������������������������������������������������������������������������������������������         ���������������         ������������������         ���������������������������������������������������������������������������������������������������������������   ���                           ���������������������������������            ������������������               ���������������                              ���������            ������         ������������                  ������������������            ������������������                           ���������������������������������                        ������            ���������������������������������               ������������������������������         ������������������������������������������������������������������������������������������������������������������������������������������         ���������������         ������������������         ���������������������������������������������������������������������������������������                           ���������������������������   ������������������������������������            ������������               ������������������������������������            ���������������������������������������������������������������������������������������������������������������������������������            ���������������������������������                     ���������            ������������      ���������������               ������������������������������         ������������������������������������������������������������������������������������������������������������������������������������������            ������������         ���������������            ���������������������������������������������������������������������������������������   ���������������������������������������������������   ������������������������������������                                    ���������������������������������������            ���������������������������������������������������������������������������������������������������������������������������������            ���������������������������������                     ���������            ������������                                 ���������������������������������         ������������������������������������������������������������������������������������������������������������������������������������������            ������������         ���������������         ������������������������������������������������������������������������������������������   ���������������������������������������������������   ������������������������������������������                           ������������������������������������������            ������������������������������������������������������������������������������������            ���������������������������������            ���������������������������������                  ������������            ������������                              ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������         ������������         ������������            ������������������������������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������                     ���������������������������������������������            ������������������������������������������������������������������������������������            ���������������������������������            ���������������������������������               ���������������            ���������������������               ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������         ���������         ���������            ���������������������������������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������������������������������������������������������������������            ������������������������������������������������������������������������������������            ���������������������������������            ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������            ���         ���               ������������������������������������������������������������������������������������������������   ���������������������������                           ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������         ���         ������         ���������������������������������������������������������������������������������������������������                           ���   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������         ������   ���������������������������������������������������������������������������������������������������������������������������������   ���   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ������������������������������������������������������������������������������������������������������������������������������������������   ���   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             ���������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���������������������         ���         ������         ������   ������         ���         ������         ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ������������������������   ���������   ���������   ���   ������   ���������   ������������   ������   ���   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ������������������������   ������������   ������   ���   ���������   ������   ������         ������   ���   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���������������������      ������         ���   ������   ���������   ���      ������   ���������   ������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ������������������������������������������������������������������   ������������������������������������������������������������������������������������������            ���            ���         ���������            ���   ���         ������������������������������������������������������������                        ���            ���������         ���   ���            ������������������������������������������������������������   ������   ���            ���   ���������   ���         ���������         ���   ���         ���������������������������������������������         ���      ���   ���   ���               ������   ���                  ���      ���������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������   ������   ���������      ���   ���   ���������������      ������      ���   ������������������������������������������������������������   ������   ���������   ���   ������   ���������������   ���������   ������   ������������������������������������������������������������   ������   ���   ������   ���   ���         ������   ���������������      ���������   ���      ������������������������������������������   ���������   ������   ���   ���               ������   ���                  ���   ������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������         ������            ���������������������������������������������������������������������������������   ������   ���         ������         ������������      ���������      ���   ������������������������������������������������������������   ������   ���      ������            ������������      ���������   ������   ������������������������������������������������������������            ���   ������   ���         ���   ������   ������������������   ���������   ���      ������������������������������������������         ���      ���         ���   ���   ���                     ���                  ���������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������   ������   ���   ������������������������������������������������������������������������������������������   ������   ���            ���   ���   ���������   ���      ���������   ���   ������������������������������������������������������������   ������   ���   ���   ���            ���������         ���������         ���������������������������������������������������������������   ������   ���            ���      ������   ������   ������������         ���������         ���������������������������������������������         ���   ������   ���������������������������������������������������������   ������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������   ������   ���   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������   ���      ���      ���   ���������������������������������������������������������������                                                                                                                     ���������������������                                                                                                                  ���������������������������                                                                                                                              ���                                                                                                                                       ���������������������������   ���������������������������������������������������   ���������������������������������������������������      ���������������   ������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ���������������������������   ������������������������������������������������������������������������������������������������������������������������   ���   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������   ���������������������������������������������������   ������������������������������������������������������������                  ���������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ���������������������������   ������������������������������������������������������������������������������������������������������������������������   ���   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������   ���������������������������������������������������   ���������������������������������������������������         ������������������      ���������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ���������������������������   ������������������������������������������������������������������������������������������������������������������������   ���   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������   ���������������������������������������������������   ���������������������������������������������      ���������������������������������      ���������������������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ���������������������������   ������������������������������������������������������������������������������������������������������������������������   ���   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������   ���������������������������������������������������   ���������������������������������������      ���������������������������������������������   ������������������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ���������������������������   ������������������������������������������������������������������������������������������������������������������������   ���   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������   ���������������������������������������������������   ������������������������������������   ������������������������������������������������������   ���������������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ���������������������������   ������������������������������������������������������������������������������������������������������������������������   ���   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������   ���������������������������������������������������   ������������������������������������   ���������������������������������������������������������   ������������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ���������������������������   ������������������������������������������������������������������������������������������������������������������������   ���   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������   ���������������������������������������������������   ���������������������������������   ������������������������������������������������������������   ������������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ���������������������������   ������������������������������������������������������������������������������������������������������������������������   ���   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������   ���������������������������������������������������   ������������������������������   ������������������������������������������������������������������   ���������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ���������������������������   ������������������������������������������������������������������������������������������������������������������������   ���   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������   ���������������������������������������������������   ������������������������������   ������������������������������������������������������������������   ���������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ���������������������������   ������������������������������������������������������������������������������������������������������������������������   ���   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������   ���������������������������                           ������������������������������   ������������������������������������������������������������������   ���������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ���������������������������   ������������������������������������������������������������������������������������������������������������������������   ���   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������                           ���   ���������������������������������������������������   ������������������������������������������������������������������������   ������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ���������������������������   ������������������������������������������������������������������������������������������������������������������������   ���   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���   ���������������������������������������������������   ������������������������������������������������������������������������   ������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ���������������������������   ������������������������������������������������������������������������������������������������������������������������   ���   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���   ���������������������������������������������������   ������������������������������������������������������������������������   ������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ���������������������������   ������������������������������������������������������������������������������������������������������������������������   ���   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���   ������������������������������������������������������   ������������������������������������������������������������������   ���������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ���������������������������   ������������������������������������������������������������������������������������������������������������������������   ���   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���   ������������������������������������������������������   ������������������������������������������������������������������   ���������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ���������������������������                                                                                                                              ���   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���   ������������������������������������������������������   ���������������������������������������������������������������   ������������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���                           ���������������������������������   ������������������������������������������������������������   ������������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������                           ���������������������������   ������������������������������������   ������������������������������������������������������   ���������������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������   ���������������������������������������������������   ������������������������������������   ������������������������������������������������������   ���������������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������   ���������������������������������������������������   ���������������������������������������   ������������������������������������������������   ������������������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������   ���������������������������������������������������   ������������������������������������������         ������������������������������         ���������������������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������   ���������������������������������������������������   ���������������������������������������������������         ������������         ������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������   ���������������������������������������������������   ������������������������������������������������������������            ���������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������   ���������������������������                           ���������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������                           ���   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���                           ���������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������                           ���������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������   ���������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                       ���������������������������   ���������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������                           ���������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                     ���������������������                                                                                                                  ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                           ���   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                            ������������������������������������������������������������������  ���   ������  ���   ������������������������������������������������������������������������������������������ �  ���   ������  ���   �?����������������������������������������������������������������������������������������������������?��������?����������w�����������w��������������������������w��������������� ������������w�������������?���������������w��������������������������{�����������{����������������{�����������{����������������w�����������{��������������{�����������{������� ��������w�����������{�����?��������{����������������������������{����������������������������w�����������{���������������{�������������w���������������{�����������{�����������������{�����������{����������� ���{��������������w���������?�����{�����������{�����������������{�����������{���������������{�����������{�������������������?���������?������������������������������������� ����������������������������?��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                            �����������������������������߿����������������������������߿�                            ������������������������������������������������������������������������������������������������������������������������������                            �����������������������������߿�                            ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                              ?���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                              �������������������������������������������������������������������������������������������������������������������������������������������������������������                            ��������������������������������������������������������������                            �����������������������������������������������������������������������������������������������                            ��������������������������������������������������������������                            ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������ ��������������������������������������������������������������������?��������?����������������������w������������������w�����������w����������������w�����������w���������������w�����������{����������� ������������������w����������������w�����������{����������������{��������������w���������������{��������������w�����������������w�����������w�����������������{������������������������������w�����������w������ ����������w�����������w����������������{�����������{������������������������������w����������������{�����������{����������������{��������������w�������������{��������������w�� �������������{���������������������?�����������������������������������������������������������������������������������������������������������������������������������������������   ���  ������   ?���  � ������������������������������������������������������������������������������������������   ���  ������   ?���  �����������������������������������                            �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                             ������������������������������������������������������������������������������������������������������������������������������������������������������������������������_�����������������������������'�_�����������������������������%�O����������������������������M��������������������o�������������������������������o����������  �      ������������������������������������������������������������������������    �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      �����������������������������������������������?���  ���������������������� ����������������������������������������������������������������������������������������������������������������������������������������������������    ������������������������������������?����������������������������� ���������������������������������������������������������������������?�>?�~ ����������������� > ?� ?�| ���������������  ?� ?�| ���������������<?<?�x���������������?�~>?�<?�x�������������� ���>>�<?�p���������?���������>?�<?�p�~ �����?���������>?<?�`�> ������?��������<?�b�> ������?��������?�B���������~?�������~ � ?���������|~?�����?�~�1�~�?���������|~?��� ���<������?�|�������<|?������� ?������?� ?�������<|������� �����?� �������<x��������������?�>���������p���������������?�������������A������?������������������������c���� ��������������������������o���������������������������������������������������������������������������������������������������������������������������������������������������������������������                               ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                             ������������������������������������������������������������������������������������������������������c�������������������������������k������������������������������lk������������������������������M�������������������������������������8������?��Ph�����������ܯ���u�����j7Ο��Ph����������я9��L<����h��������������Ю���T8����	��?�����������������������������������������/���    �    �     �    ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������?����������������������������� ���������������������������������������������������������������������������������������������������������������������������������������������������     �����������������������������������������?����������������������������� ������������������������������������������������������������������������������������������������������������������������������������������������������������������?����������������������������?����������������������������� �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������?����������������������������� ���������������������������������������������������������    ���������������������������������������������������������������������������������������������������?������    �    ������������� �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                               ��������������������������������NNNNN                                                                                                                             Cadlink Version 6.1
 �P�B��+E�L̞3��$h��Uq��
�!M[�r�I0?�쪙O˻=���W1r��Q�=����|�8YZ0��Y�D��v�v���f�2dz�%&�-��_yy%'P�n�!A��I�f�&P°)C�N <   �G��b�����޲ ŷ�a�<��� po������x�g��}KCU�p������g ��I�3�9������'Pzp�7�<HB'<�?����fN1lʀ���4=�d\i.�9�_P�n�����>���}�C�}@˯ x��Cؔ	#��8��w��$�3�Y���Or�f�?af�ZHr2|zNF�z82"gR��0g2wB��83�qfR�,�9Y��Do� 9�3��"�#�>��$!�9eʸ�&'¦wAN����!'�9�$gl?�8��a���]hCZHs(���)�!3|CfHr;�d?N)�C�:e���u�D�x8�2"�2'B�#pg���?��9S���ІĐ�PD�����G��LC�qmȌ|�d�y<�02ef�$d�13�q?!̎�	����x"'��3e�
�a�=D8���ƈ�
e�
G���ǩ��!��  )1��ឆ �=�2e��J���^�~��{4�����'7q�I�3sLs/F���=3A�%��_r�� ½z�Ls/F���=MA�{�fL���_pឬ �=g̘�`��^�~��{̂�hʔ�Cv`�{1��"�ӌ�܁i���\�0�p���܋�/�pc��p���܋�/�pOf�3sLs/F���=�A�{�1c��<0ͽ�����9c����4�b�.��D�W�i���\��9�p��L�?����_p�� �=3f���^�~��{̃�4c��{`�{1��"�sƌ��i���$������^����K$�����_ �{��/D��2� ��P�/$����
�� �1�
��]S�	ua�?D�����h�p�r��_Hr�g���?����I��B��a�"D8�S�@a�@��Ot��Ay����׹7?!����@��	B�M7kK�0l��y����СS O�
�(V@���b�1l���5`��&yhY/0`�eZ���躻�#g�Ls�Y�b����ֽ���2o�%�Tmr{F�0�z�-<!R�L͈Q�� @ l �pv6o��?r �`@ٿM�z��a` �oF �0����uD �n �,�XS � �&�@v��5��o�]�M��	A��С	��D��� �d��r��YyP hk� ���� ��c{V � ���$��{@�	�;$�2ʗ{<${�c��s:���(�T��K��?2��ɔO��n�]�?����?�#��� ׃�C � �@ s � �kkM ��Vnp����_��8: �޵yL�y�f�}m��uG )}2�*;���vV;;���#v��bhЏ�,�!����!�0`zc�0q�	�DF����{�����/�,@�0P��¸ po��~!|�/^�;r��'B�4P+�D���4��7DJ��*/�?��s��#T�U���<4e��!�O���͟��Wr�^3f�0�|����'��̘��<<�G�Ռ����|�M~F:D�0dN�Pa
<%�Ѓ��{� <qb$)�#A��@����i$�O��SWFF���}L�Pq�S�La�ԟ!N�P͇J(Lc��7#�0j6�4\�GC�.�S�4b�p�vTJ0%C��!y"Di����F��U 3��P���Y��Z?�1b�O(T�6�nZs8j=�g"CMo��9�0:�Q9j<� �	�CO�� ���#|���DG��PA:�%W�m��5`Ġq�F��oh��Q��8	X�jݶӫ��Z}3�h0\��k�Ō2�
���QCf���M���B�����Z���@9rܰ��a}R�Q���2T#g{l䤅l̸1g�7��nм�8j�ҍ�U^�~�rẬ�:�k������]4f�a��l@L)\P�<����cb�gǸ�k����6i��e������r�S�Y�5���ې����唳��;6���]X���F9���X���#��T�ŵ~��]�dԐI8�L�,N5���L�f̘����Ζ_?9dѺ��Jo�+�cy,`[/�U�{	Io���4��䐳����j�K�������o���,�n.�i��Wv�Y9��f�bF������2RS+!y"D��X��}q�ل"P�HiZ�dH��[e&,X��D����N���_L�����jA=�,666z�&
�thTn�F�も��2���Q��^ך��pN獡�ל�F��4����.�ްhN�)b��'�AQ��^��f`6:��o\F�)
u����F̘b�n��f���1�Ɛ���|4c��v�$ܰ�M�PW�cn��7��(�E����A�����xM�YKDbи	����pj�,F�ᲘC�.�o��7nРٸ�(p��ͺ���ҎLTX8��ܕ�uA�2z�'���%�����ƀ�׍�ï1m2p��B5+Z�o��T'z!�ܰ�������!QgFN��0�l#��/����'8nĄÿ��S���6����1���	g��\Y6l�D栖(օ@]t����]���W'D
����P(��و��BaTRG�5��q���74*#�	�'B�X�V�۠�*M�Pi�-17d��qd�aF��)���	��dF� 9τI*N������i{1��d
���TIB���^=���<�W��גY�Ȍ�n��7pVȘf[9s��3�^���T^޵�s.pg�x�Q���d��'c�6l�~�W30�&rȌ�p��1S��pY��omȠY�h����
F#G��,`�o��f�O�z��:ɷ#�~�Y]2<�\���g�V�F�m��lr�6�6 �&���³���7SuX%3�kf	�q2�z/f8b�7�Q���8�Ζ�+x�Ŭ�+"f
͸q�eԿ[jz�ĺ��z�Y�h�peWj����1�&�d�y�]�Z��c���ʮ�=O�fݖ¹lf9l��Y�ͻ!s��2��f��\pV�lh�М�봹�9�ֺV6N�Gh�ӆ�	�h�#:nՄa�D"�3\�׷U��c��\�l�n����h!Ez�p̐�V�ר��5�#�8�*'^��!Z'4�B^�E`��Y�ḧ4T�i�6�f�lĠ)v�L+ՄD)������Z�*�9	�1cM�:���"6j�	uu��3c��gi�aӮ����as$YՕ(�G9���`���;ɘ)�0�л�G��B�2>����e�n��Jn����@k�@N$5�p�c�_�1�3lڥ����Ā�CftS]��qv��\8��lۄ9f̬MX
�Ԏ�}�׺0L��+���]3!Q&7�:5���:3r*(�Y�6����/���1m�!�B�NN�o�lа!C&���L��U���.�PTҒֱ1C��'�u��lਉ�J���D���EU'�[[F&D
�r*��!P�T}� p}�ۉY&h����׭�TF.<�D�p<)݄�����p�ƌ���{��>�/p��\�B�S�8�N�$O�(Yb`��=0r6�J� To]:@&�.l�t,4\6�n�*R@F�9����H�F1�B�iRc�T?S�<m/f{C�L=���TIB���^=���?r�R��.0�79r�,�%�.���Ɗ���]V7��(eZ"���-��xas��Fa�Vp���A5�Z"�Ȍ���&Ե<W�T�Cf4f�@�,����%�7�mRG,��]o6pV3	c�ȩ2�7J��Yغ��5PC&<�jĀ_�䬓31Z/s6K��(4$��Cfܘ	J�����A��w�47S5��ńIs0U�=�e8�V�I9E��y���|����2`�E��0R�4��8�ńC�w�i/&<ơ�S!Lj��S#F8��j�c&^9�1ZGC�B]�(�r]Ō*l��,��9���dF5b��i-؄���+�-�S+&N�qTdÆ�3�
��x�ȰAcȍ 7n��S.f�E7T���d�D-$3���`�,	8f"˽pL��!�	S%��I���:�Y6n"h�En�R���pk�l¯�:�	���A�S}9�q��"�!Bp�=0AH�M��QA��p��)41j�q�9|Մ�N�ƨ���72f 9�*	RG�.EA�ZbB�Z`B�Zf�O�uBj�a�Zo�0�0&�0n�"��`fq���t�lR7��7#�b�^3�t�6��Z- d��a��(ޠ���a�;6p�B�8��Y@�M�32�,��P�:
W��(3�7j��	�םM�����X��%g�����j�T�4�]11��3���x��ݐD��	y�'��{�ɴ+o�Sbܸ3(.�tTc�쟮��[�ɼ�&�L�Y����D�/r]��e��W�1��!8f�J�0A@�Ԑm)1�4K��1f"iY��4�Ĝ�l�K������k��zm����1�N��"|h���}9��F�D�44�j8pȠ1#'C~D���UڠQ�f��Ũ��� 5�!R$'i��!�MX34j1S��Cf�h��j��f��9E��k��i��hB]�mհ�ʁc�`���1JM4�"�����X̦�2�P���xY�a#2rⵕ�!A`!
}m�4�/�d�,)6`��B�˲E�F�R:��,2���B9/�
�=8j����q�
MŬ� ���f
83��L����NN���԰IjG̺mb}��k�h,)8���<,FrE˒�3�/J5j6�&k��h���!����2�3�"fTx���q��0U�5��Fݬ}�Řacf�r���xU	���#$(�P��'�KUY'5�y�ЄYf2S�&��U�ͭ���G�*d1�!1!�
��T[�n�����»4�40�q#W\	��C̂"fAY8C��L��E~3l��3�R�g1\�܄�uGn�&��MXꢋE���.nDv(jat��}3a�<RaTg�,L��M�q���	�#����r*L�a@F�@!R�/��ʈ>C�D��3ʍ3pب�<*M��k�@D��:1����E̚�BEj�`�aHA���l�,T�&5&N�3����/7���SoJ�$D��^=�4��!��GL�g���r_�`�,����#G͞�}9n��[���R��4[�Y ܈q����1]�m*шӕ��'<��M��fl����L�c=7�&^%A��#H��PW)�+�5�ܭwcnĄ���c4G4k�&r�y�������
1#&L�hF�����:o�LR{6��w���2b��	>�3�"G�<�ך�Z1qԊ�ط�C��R&Nx�$�ҦO8˖M�J�\�r|Tb�ѷ�p3T[w3�5l�Ȅ�죂������ud���X�#P�!D�� R$&8iϦj����5�&<�˩�/lkhf��R�j��0q3¢�:�)گ�e*&��dȬ�
Yu1h.��+��Q0Ҝ2Us7�!#&������77\M84_w4Us6d̸Q���O5�S5Ws=�dV�ᬼ5fVKN��b̬ 5�� 
N���.mg�ʴ�\	��g��52�YU�{u�)2�;�*��ٴ8nb4g����{7�����͗���حF�m^nj����ƂuA�`����`�ٌp^��93�)t3B��j6�`�P�̆.���X�*k �"7n�U��*l­J��	�*����f ��ܐ��d�DP��J��|�p3�Cj��������0���s1cFM�[{DfV�Q�Q�͒2ÅL�*l J��	*�	*�	�*rؠ��4�īAh�2�F� ���P�M��X4aWcԄA4l^sW�U@Dh񒁳TX�ڕ������f�iA�d�L�9`ܘY:	�P��%�e4�����(��o�\�8h̸��&5VO�CK�Lȫp 'S�`��lá}��pN�f�٬���Da�47���1�FL�#�!9bB]��LK�͹��4�1n���Wu!J٢;uS�Gf}�	c�B��\�D���"c�U�.^+4+/H�"6�B_�ԅm51���bsG�(��s�'� ��EѨ����1cfCd�l��x��0R��9p��F�WZ�+���O���$-a`V�v�؄�.�US2`V���p%�Т������4�� G�m�X8����gѡ9�#�"rU�l�rĜ`+��D�FD���P�L��`7r��r��6�ͣY�0hبa#���n��b�<�bx�8r�n���j�R��jЬ�f�P�"��&`�r_����7�F�r��kn�"D�����ҜL4�eS�^�w��=A��}����uj�֡��[3�7h"Թ	K]�i����+�͖j��@�N�b
�̰9D.��Zљ���-��b��=s�P*�b��0�)��*�"zt�"q �cQ#;�$�p(ZaDg�,L��M�qC���08�.�	NFt-eT��� �P�DH�Q��j���#���*M�P0���4��ׄ���W�Y��T
�̓���S_�5�6��*L�	   ��?�������^�e�o��@yu�/ �� ���#|�D���#I���@1!T���O�j�x¯&Y�8�0q��)L��?E4a��	0�0���� uRb�)��c*�pq��3h�c��:ۃW9��ƌ3p�l5/�����1jĬ�A\�����f7�93k$�U,0�Ed��o8#��z�b�f�0h޴	�H:t�b�p޹{�X%.O��6+��̚����,�M�acf�o%G���W��n�'�8\ܬ�ƶ����7k'��L�o���Ͱ�7d6��l��X�*`V#�Ο�N=�u�|{%��ey��p��Y���r�l7{Ĭ�:��M�Ynʕ��r�ؾ3��x6a抨Y�Zղ���e�fuW����Xw2b�,��2b�Yz+��WT��;z_�D�p��]#0Q�o��^fj��f��n.��Y�etxɺ.E8l�m+8�oɳ�ݭ��z�YM9+�&������7eAZ��7nn�&��{�	�j��mxY�Y��F�Y>j^�̸�"f�et��b��b�"�L\�SFF�bهs��ѫs����n�j�Zb������@ѱ��P1xXl~��˚Mt����s�y@0�ck|q5�Q��+ھi\��=ǖ�p��?�2��Yo3l�,���T�%ZOj��5?5<8'�r٠�<V���,�[M��$�P\��ՠCtž�u]0�'�e�D���4l��٣��@�w)-�j��fج���d�u?���y�Kt�����=��'�>�����Qs���q���R�ES���̄��P�!���|��$'���\2�-��a�e;1r�2�<��(Ʈ���ńf���c�����g��[l&:�7���/��-Ѩ	�����h2���f�
�r�Y��-͒$��Fs���R!�tV��d�^٥���i�����N1\n��5uszcxعZ�IΠy������C����j�_��m�Ya`V�2�沨BU's�5��_�f��,��~��_2����`�<���łf1>�Pi�
H�r�[�ᰑ3 ������+�������B���(&Y�8MzL��g
����7C�L=���V�����T.n��~XX�uZp�h�/r6%g�t�_�
t�F�&��}�C�L$�]E��b
#*ȇ1b,KrN1E���J4oڄ	`��\�ы���3����چ̚����	hذ1�ܷ������a�x�G@R�_.���Ɂ�<������>0hܐAl�Y0��Pg@/�S�6�^�!�fYެ5\�f� �Jn��f�_�{�	2K��B��۽SN$�s@>�m��Q'��4֝�6�z����m���-�U#��W9�9����D"W�EW3�K7���2:�d]�"6϶�˷�� ��Vnj�ᬦ��k$}Wa�oʂ�f�/2n���M���"�!����Bp��D6���Q�6`ƽ1.�#���Qe�
�22r�>��U�^�c���EpSW���D�������ğ�����`��t]�l��u����	[㋫ɏZM^���H�P��9�$���M�q��Y���z�a�f��f�-�zR�Ĭ�����9Q��������fQ_�j�$&iP��j�ͭ�+�լ낱<�,�%"'e��Рa���5��� ��Ki!U�T7�f���(�'���q.G��\��;����<�8���}W�ό�3,�؎+��ސj,��m4d&��4��X7'9�E��:��nI�.ۉ������D1v�6�P.&4��fh��7��>���b3ѱ��Mm~?m�FM�̎P\�F��~�6;W �C̺/n9h�$�l6�C��
���j ��.�u_HN�M$v��r�嬩�C����պOr���T���x���nW���"]n�
�B��4�E*X�:������r�7��f����f��Q�������'�7��&Pi�
H�r�βe��7p_�z+��������H"1�0L�Pq�8�8��&O۟��8�z��A=w��$�Bs��As.�W~#�ɭ��F؈�� �13@��nt�h�1K��H������T�c�X�b�F�0h޴	�H:t�b�ȯ3y5��a��J樓��.�nV4�2�ܷ�����	a�x�G@Z�_.���Ɂ�M�S��a�4nν���*`V#�΀fT�*��R{u���j��5��j2�-�[����\_7jVh�1d�l�pt��a`i��M��f��Y��&g5��9�D���ZQ\nк!�X6p��� w�fv׃LX�����F�}2lB��Kφ���o�C���&�Y�Ճ�F�9r6u������lR6��&��%af�[x��=�/�s��39��Ɩ ͆W~!����&��rؼf�����l�&���p�M6�L��@,k8�5����䍭!���fᔃ��I�	7\����d�7*&�<.��zWj�#�������� k�h�er��b��b��
.��s!Y����N6����P������B�&���J�D�I$��j�a�`��b���l`=W��n窲Q�1Ic"Wc�dUS�<����&#�M6��v/�l�.��sT�+�c{Qm��b�D2~;.d�L6�V)�`.j�{r�16�Y���ktt�Y&acC��j�0�d4l*�L(8�
2�kON��&��٬��Ӆ̒Y�`�,�Ua�Hf���v��b]��f3�3[.hVa����G稙Mm^��_�-�,�p����}���p*GW ���Ž��$��.�͛���Y55��Y��XN�M$Ί�"g�9<.��s�j������'a��z�V`�Dgg|���3���X8:�x��Y�K��ˡ
,T���@�dm���������W������M<�%_y2�@�I* �����!E�P��L=�"D�-��b���Ӵc�T?S�<m��d�	����$L�n�lN����>~�����l7�.0��a9/_ 7�f��w���#��*<S��o8#Ʋ �S4�X��A�M� F�С�����ud��:8WF���e��;6af�[�Qfe���0{;�# ��/�f���A�&Ϳ).?�s`A��Y0��Pe@'�S�ȩ^�YH���������-p�ui-�n��YO1��M�9�۞����K��s��e\ r�19l��y�U��jVv�� ]C3�6\`�������.s6��_8��e�<�1�ѲpbA�~髑#f�i��mV�b]ak��Qv�Հsk7��@�<	3f�x#`ntJ�岎r�٬<�e"'��K�"F�fW��	S�D-�F�A���z|��\�y�9���Z_2`�,XK�̧E�` 9j���.�Ű��.��Ņ��O�~��5r�вb6,�{օP�Ȧ����V��'������䛒M� ���pY ��3�����|K�,e2��v'����y��f�x�o����V9`�@5f����as��Y!��f�F_˵&s8X/3эE�^O��w�a38�8-&�de�)�7�aP�7)&��ͺ�Y���Yr�D1x���b�&��%L^�e�v0�Rѱ lX���`/e�0�{g.��*ͦ7�H�ę,���s��, A{b�{�]m.����7��l*6.�a��7k����.�
����14+���f��y��FL�ݸy��U_9�\�1|p<ŏ��b���\Ȭ��X����|F#�]X�4�pYH�n��r��F�P�B���Y��H��_��y��SV��MXH�Q���7���&A��d���Y��9I�� �a��*��������e,H!4�6�I*N�����i���d�1����$�m�I��!�,4n.ĕ\���s�ɬ����a�̦���lt�h�31`���*\�Z&�cY�jY4�X��A�M� F�С�ﾂ�Nv4l�z��6��.ˎ�r3�Q6f��Vr�Yپ -�Ǉ�c��PM�P$��r1n�8hФ�7�e�f�l	�Ӡ��)1���B.�v9)�,�3�2-bY"�Z��W�l��0��/}7)0l�f���D7�fa[N������&�9�?�кF��Z:���p�Y��E.'�L�e��u�c�$G����|��
�lRC�TC��e��T��Np���Ʈ�];��� �9ϸ��Wwz�Ѩ9�F0w�����܂��
��M�1cF���Zڛ�FMJ�Se��i��Y��r�&��d��YrlЬ�ټ���_\�vS�^��+�M�H1ۑY,� �l���>1��DX��̉��<к�٘����Z���F�,�yɸ��d�٨H	�'&��H���p�]���YP��Q7]ϵ^ߵR������hˢ}�' �"��]����X\�l��&3a��kVd�?p<8�%��S{m���wєI���FNdͬ⊯��7m��Y�%��:�9�6GLD��Ԭ�]9G78��	�#W�܈j����|��Ǥ�0�����W����ޟ@p�תnsB��\O��BG��T�a�L�ؽc�fF�܌��&��W��o=�I�@5Bq5Y�b26��˒Y���\1��C���9�T6~`Y�+��I�)�Q5�L�|	P��ʺY�巾l̠�l��_�%�!3�+F��p����|s
��T,�Y�� ft?l���MfÅ�1t���`.( j�p9��ٺ�9f�(֮�ca��kM�qjY�˷���[jn���9���j�{�;5`���f�؄$�D-.�s&a�^P �1��e��P-/2fV�L0�^�̄�d6��m\���u^4\Vw���P��A�U^5�ҳ��J.lG�
���I��-{2� .�28���x01��'�m9?��&G�B �L!���p�M\�0�M��l�n�z���7T*X�:��6�B�gAY���a�ϻ�������_M��gH�Q�1h��l�&A��Ĺ�*Rۃ���p���BR/$C�c����b�T?S�<m�q2��ۃR�L"BuLB2����p�Dg�;66�f�pof �m�f}ќ!��?�U$x*�0��F�eA�)��2�P	��M�0���C�+����ްJp��8d��!��1�pY.d6g�^��V9ʬl_�f�'����9`��5"SP��F6 ����mH�r`�8l�ȣc]��U[�԰��X37rڳ�a	%h��C7jR0C�yo�Al�,�;.gK��h�53��_�n����^��uŖ��kh��%�	2r`EG4�Y�z�02`Ј�kn^��e����������E�@*��Rק�|C�����,¥tC�f7�:�ͦWwo,��p�U�]�~�l��-�L�94Ϸ��	��{Zn��.����𫴦f���I�m��/���Q���0~/Z6\��e��7�R�4�,}1�{����l�.���?owݐ���������>�Kj<0\�ꍽqy�6���&\FDq�q�b*+�sa}�v�Z�l�`Cf�Ѣ9����bf1�us*�M4n��r6�n�}Z�I���\���Iu8���Qs�\����
0�%3\�Q�j.ǡi�X[����CM��e��B�f�9E�"Z�%w�������"��uwk	l820�Y�r�lȜEIV,8��@vv�قG&:�\8dVY��]'1acA|qƈ��*%�3u�N���Lp3d*����L�3TM

?�,��9{ΕE�FL$"�h�Ԓ�Y�b��15g�v[�	K�jo#h��b��8��Wcnf5�B_�9���
�8Dc&��X8�,�M/��9����ڭ��;4�h��}�p������#���ۨ��X�f�acG|q5{(�f�)X�;���K��6�هZ4N2��֫q��8��y�3r�Dc�"Y��l=��e;p����K���f��l��覣�e�W_ͺ�D�p�����t5�����~.�5�˵P����Y���No�8�[4/\��t��L��]W2��i�����0nj�h�$�63y7����첉nt�a3:��m� �yFf �B���\U�`��d� ��l��ٿy��Uޫ� }kb��$O�(��BVnE��T������fb��	F�%Sg=�BEj}���_zK��s�zN2d�l�I*N�����i�s�'S��=(53Xn�&��^�nɘ��ݤ.#��&��/���Q�u?��$�ey��.k�f��;� 	v	�)���c�x��|E���J4oڄ	`��\�����w�䰹b`V���pYvd���U��eVBqa�x������:��9Ք��b�<�9�����Y�d����.1�f5����Ti6j*H�Q��LN5�r�&��iu,��]ACf�;x9ܯ�z�q�Jf�Ң�nE��Bղǜ5C���b����I�Y0+dWNdD�!\ ����V_x��1f����[g8/H�RΪ����n�pY�ŰKt���P0zb,�9#�U^Q3��>$m�"nd�ň�6�㋫�7�������%Nx���{��3�}��T$�#�h�֓ts�F�%[Vl�Dd�V�82E1HLҠ�ՠ�[:����}����^n̼��#dn�8d�,���,93@؜pr�,55��䎔(���VU�)Z��C�һU爘Lf���4���jy�����D6|)�lw�l�Ś���1*���l��=�Ư.���?��Et�l����d�f�D2\���4�krԌ�lVvC+�z/�p���lI�U7`���e�esn�{e��������l����
��&�;|F�i=����D_��4g��x��fQɑ#g�p�lDL$�v�3����{c��3S��k�d��eA�sIN�=��|��Q�.����\����~9Ku�T����ӝ�@�h�k�OfS�`��G�?a y"D�3�K��ωJ� T@R�B5��"�,4G���R
�����+H�EL�Pq��8��&O��C�L=���V�L�����V��"�^�a���Yvd���ђ6�F��р9�}j�f~q�]E�wb
�+��1b,�s�̘��J4oڄ	`��\�Q3��}�U�B�	-ƍ�C�lvّ9��a�f#j���������x�GA}�/_�k'4i~1Xf�l	�2��E1��$L�&�S��i������N����k�`����3����f���z�u�Y�.���d\��(�!�faX�M����#9�c��,{7K~�f������`)����g�f9�7�d�~�Ԅ�#W�Ԫ��^ʑs��������F�u^��q7_߸�-�1��{#���É?A,1kof�f�<��3sբ�!@�L��u�|s�,P7%5��BUt @�,��ٟ(�<�t����Zo�&A�\@�t��N��|Ѩ�Bf!}E�P�Z0���F�"0�6�QN�$a�N    4���'�w��އ������{b� |���>L�Pq1q��)L��?qQA2�j>W���>M�$ij�M)(R�j��K�N�\uP�ֹ��U��oGH-I@�_��Q�����0l؀�c�L=� F����qsh���3`Q j����f���sp�˱^��4fb����I����{ő�nN���Z�����t��Σ�ѲЮ7�Ԗ_�k���[���{�^H��T��ā����%)�*�ً�Y����Emq�$�Lj��W�?7���l^��dCfᒓ`�&��^�l0��hR%'�Z/�N5�g�&.�%��x�X/1p����TA��2b�lRM��b^gq����Y���0g�[�,5bR%ǅ�
&Ů�W�Y7`<2s�,2Y=�D�(������bUCƍ�9�D� se��sn�$,��:�H�!����ؠ��r)FQZ�p=J��4g�+̀9H&���v�S,^c1�PME�V3q��9��$8���L��H�_�h#���o��u��YVp�8H(��MFܬ�d�z=%3)T�����+NF�u��q��,91a٠A�FN������2k+MI���k!_�6df�CN�u��M�3���e2W���f�6Hf e)�
�h@�4�d��Ĝ*k�: `���%�&�gh�f���K�"�\3��4b��� cf�j"P-�u��91�8;1��1sR�f�ꫲx2�żd��$��9l��@89\���BX��%rXJ�T���J!n tlB'�D���q� ��J���xܰI���F�&��(ÚC��Ȣ��N�V}$Rn����J���%�FN�I�q�y�A7��I��⠲�T��$N��ZW+�6��,59)������\	0h��Iv�1���ӲZ���ƊIj"g�c&D�H���W�9�.��D�*2�����h�m��Y�B͐���0��P�jԘ�q(3�᫋Xqr�Y7fҎ6�e��"P}1�.�------------===== CDL4 =====BM�      �   |                                 �  �  �        niW0L�г� a� �.nd]��z �Ը ��I �O�                        ������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         ���������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������   ���������������������������                                                                                       ������������������������������������������������������������������������                                                                              ���������������������������������������������������������������������������������������������������������������������������������������������������                                                                           ������������������������������������������������������������������������                                                                                          ���������������������������   ���������������������������������������������������������������������������������������   ���������������������������   ���������������������������������������������������������������������������������   ������������������������������������������������������������������������   ������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������   ������������������������������������������������������������������������   ������������������������������������������������������������������������������������   ���������������������������   ���������������������������������������������������������������������������������������   ���������������������������   ���������������������������������������������������������������������������������   ������������������������������������������������������������������������   ������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������   ������������������������������������������������������������������������   ������������������������������������������������������������������������������������   ���������������������������   ���������������������������������������������������������������������������������������   ���������������������������   ���������������������������������������������������������������������������������   ������������������������������������������������������������������������   ������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������   ������������������������������������������������������������������������   ������������������������������������������������������������������������������������   ���������������������������   ���������������������������������������������������������������                           ���������������������������                                                                                       ������������������������������������������������������������������������                                                                              ���������������������������������������������������������������������������������������������������������������������������������������������������                                                                           ������������������������������������������������������������������������                                                                                          ���������������������������                        ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ���������������������������������������������������������������������������������������������               ���������������������������                  ���������������������������                  ���������������������������                  ���������������������������                  ���������������������������                  ���������������������������               ������������������������������               ������������������������������               ������������������������������               ������������������������������               ���������������������������                  ���������������������������                  ���������������������������������������������������������������������������   ������������������������������������������   ���������������������������������������������������������������������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ������������������������������������������������������������������������������   ������������������������������������������                           ������������������������������������������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������������������������������������                        ������������������������������������������������������������������   ���������������������������������������������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������������������������������������   ���������������������������������������������������������������������������������������   ���������������������������������������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ������������������������������������������������������������   ���������������������������������������������������������������������������������������   ���������������������������������������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ������������������������������������������������������������   ���������������������������������������������������������������������������������������   ������������������������������������������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ������������������������������������������������������������   ���������������������������������������������������������������������������������������   ������������������������������������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������������������������������������������   ���������������������������������������������������������������                           ���������������������������������������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������������������������������������������                        ������������������������������������������   ���������������������������������������������������������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������������������������������������������������������������������   ������������������������������������������   ���������������������������������������������������������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ������������������������������������������������������������������������������������������   ������������������������������������������   ���������������������������������������������������������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ������������������������������������������������������������������������������������������   ������������������������������������������   ���������������������������������������������������������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ������������������������������������������������������������������������������������������   ������������������������������������������                           ���������������������������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ������������������������������������������������������������������������                        ������������������������������������������������������������������   ������������������������������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ������������������������������������������������������������������������   ���������������������������������������������������������������������������������������   ������������������������������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ������������������������������������������������������������������������   ���������������������������������������������������������������������������������������   ���������������������������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������������������������������������������������������   ���������������������������������������������������������������������������������������   ���������������������������������������������                  ���������������������������                  ���������������������������                  ���������������������������               ������������������������������               ������������������������������               ������������������������������               ���������������������������                  ���������������������������                  ���������������������������                  ���������������������������                  ���������������������������                  ���������������������������                  ���������������������������������������������������������������������������   ���������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������                           ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                        ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ���������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         ������������������   ������������������������������������������   ���������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������   ������������������������������������������   ���������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������   ������������������������������������������   ���������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         ������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ���������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         ������������������   ������������������������������������������   ���������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������   ������������������������������������������   ���������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         ������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         ���������������������   ������������������������������������������   ������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������   ������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������   ������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         ���������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         ���������������������   ������������������������������������������   ������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������   ������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������   ������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         ���������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������                        ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                           ���������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������   ������������������������������������������������               ���������������������������                  ���������������������������                  ���������������������������                  ���������������������������                  ���������������������������                  ���������������������������               ������������������������������               ������������������������������               ������������������������������               ���������������������������                  ���������������������������                  ���������������������������                  ���������������������������������������������������������������������������   ���������������������������������������������������������������������������������������   ������������������������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������������������������������������������������������   ���������������������������������������������������������������������������������������   ���������������������������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ������������������������������������������������������������������������   ���������������������������������������������������������������������������������������   ���������������������������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ������������������������������������������������������������������������   ������������������������������������������������������������������                        ���������������������������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������������������������������������������������                           ������������������������������������������   ���������������������������������������������������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������������������������������������������������������������������������   ������������������������������������������   ���������������������������������������������������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������������������������������������������������������������������   ������������������������������������������   ���������������������������������������������������������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������������������������������������������������������������������   ������������������������������������������                        ������������������������������������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������������������������������������������                           ���������������������������������������������������������������   ������������������������������������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������������������������������������������   ���������������������������������������������������������������������������������������   ���������������������������������������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ������������������������������������������������������������   ���������������������������������������������������������������������������������������   ���������������������������������������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������������������������������������   ���������������������������������������������������������������������������������������   ������������������������������������������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������������������������������������   ���������������������������������������������������������������������������������������   ������������������������������������������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������������������������������������   ������������������������������������������������������������������                        ������������������������������������������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������������������������������������                           ������������������������������������������   ������������������������������������������������������������������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ������������   ���������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������   ���������   ������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������               ������������������������������               ������������������������������               ������������������������������               ���������������������������                  ���������������������������                  ���������������������������                  ���������������������������                  ���������������������������                  ���������������������������               ������������������������������               ������������������������������               ������������������������������               ������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������                        ���������������������������                                                                                       ���������������������������������������������������������������������������                                                                           ���������������������������������������������������������������������������������������������������������������������������������������������������                                                                              ������������������������������������������������������������������������                                                                                       ���������������������������                           ���������������������������������������������������������������   ���������������������������   ���������������������������������������������������������������������������������   ���������������������������������������������������������������������������   ���������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������   ������������������������������������������������������������������������   ���������������������������������������������������������������������������������   ���������������������������   ���������������������������������������������������������������������������������������   ���������������������������   ���������������������������������������������������������������������������������   ���������������������������������������������������������������������������   ���������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������   ������������������������������������������������������������������������   ���������������������������������������������������������������������������������   ���������������������������   ���������������������������������������������������������������������������������������   ���������������������������   ���������������������������������������������������������������������������������   ���������������������������������������������������������������������������   ���������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������   ������������������������������������������������������������������������   ���������������������������������������������������������������������������������   ���������������������������   ���������������������������������������������������������������������������������������   ���������������������������                                                                                       ���������������������������������������������������������������������������                                                                           ���������������������������������������������������������������������������������������������������������������������������������������������������                                                                              ������������������������������������������������������������������������                                                                                       ���������������������������   ���������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             ���������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������������������������������������������������   ������      ���������   ������   ���         ���   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������������������������������������������         ���      ������������   ������   ���   ���   ���   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������������������������������������������         ���      ���   ���������      ������   ���   ���      ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���      ���            ���������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������������������������������������������      ���      ������   ���������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������         ���   ������   ���������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ���������   ������   ���������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������������������������������������������                                                               ������������������������������                                                                                                                                                      ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������         ���         ������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������������������������������������������   ���������������������������������������������������������   ������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������������������������������������������   ���������������������������������������������������������   ������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                      ������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������������������������������������������   ���������������������������������������������������������   ������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������������   ������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������������������������������������������   ���������������������������������������������������������   ������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������������   ������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������������������������������������������   ���������������������������������������������������������   ������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������������   ������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������������������������������������������   ���������������������������������������������������������   ������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������������   ������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������������������������������������������   ���������������������������������������������������������   ������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������������   ������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������������������������������������������   ���������������������������������������������������������   ������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������      ������������������������������������������������   ������������������������������������������������������������������������������������������������   ������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������������������������������������������   ���������������������������������������������������������   ������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������      ������      ������������������������������������������   ������������������������������������������������������������������������������������������������   ������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������������������������������������������   ���������������������������������������������������������   ������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������      ������������������      ������������������������������������   ������������������������������������������������������������������������������������������������   ������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������������������������������������������   ���������������������������������������������������������   ������������������������������                                                                                                                                                      ���������������������������������������������������������������������������������������������������������������������������������������������      ������������������������������      ������������������������������   ������������������������������������������������������������������������������������������������   ������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������������������������������������������   ���������������������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ���������������������������   ������������������������������������������������������������������������������������������������   ������������������������������������������������������������������   ���������������������������                           ���������������������������������������������������������������������������������������                                                               ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������������   ������������������������   ������������������������������������������������������������������������������������������������   ������������������������������������������������������������������                           ���   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ������������������������   ������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������   ���   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������   ���   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������   ���   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������   ���   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������������������   ���������������������                                                                                                      ������������������������������������������������������������������������������������������   ���   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���                           ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                           ���������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������                     ������������������������               ������            ���������            ������������������������                        ���������������            ���������������               ���            ���������������������������������            ������������������            ������������                                       ���������������������������������������������������������������������������������   ���������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ������������������������������������                                    ���������������                                    ���������            ���������������������                              ������������            ������������                                 ���������������������������������            ���������������               ������������                                       ���������������������������         ������������������������������������������������   ���������������������������������   ���������������������������������������������������������������������                        ���������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ������������������������������������                                       ������������                                    ���������            ���������������������                                 ���������            ������������                                 ���������������������������������            ���������������               ������������                                       ���������������������������         ���������������������������������������������������            ���������            ���������������������������������������������������������������������                                 ���������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������               ������������                  ������               ������������            ���������            ������������������            ������������            ���������            ���������            ������������            ���������������������������������            ������������                  ���������������               ������������������������������������������������         ���������������������������������������������������������������         ���������������������������������������������������������������������������                                          ������������������������������������������������������������������������������������������������   ���������������������������                           ������������������������������               ������������������               ������            ���������������            ���������            ������������������            ���������������            ������            ���������            ������������            ���������������������������������            ������������                  ���������������������               ������������������������������������������         ������������������������������������������������������������������������������������������������������������������������������������������������            ������������������������            ���������������������������������������������������������������������������������������������                           ���   ������������������������������������������������������               ���������������������               ���            ���������������            ���������            ���������������               ���������������            ������            ������               ������������            ���������������������������������            ���������                     ������������������������               ���������������������������������������         ���������������������������������������������������������������������������������������������������������������������������������������������         ���������������������������������            ������������������������������������������������������������������������������������������������������������������   ���   ������������������������������������������������������            ������������������������               ���            ���������������            ���������            ������������������            ���������������            ������            ������               ������������            ���������������������������������            ���������                     ���������������������������               ������������������                                             ������������������������������������������������������������������������������������������������������������������������            ������������������������������������         ������������������������������������������������������������������������������������������������������������������   ���   ������������������������������������������������������            ������������������������               ���            ���������������            ���������            ������������������            ������������               ������            ������               ������������            ���������������������������������            ������                        ������������������������������               ���������������                                             ������������������������������������������������������������������������������������������������������������������������         ���������������������������������������            ���������������������������������������������������������������������������������������������������������������   ���   ������������������������������������������������������            ������������������������               ���               ������������            ���������               ���������������            ������������            ���������            ���������            ������������            ���������������������������������            ������         ���            ���������������������������������            ���������������                                             ������������������������������������������������������������������������������������������������������������������������         ������������������������������������������         ���������������������������������������������������������������������������������������������������������������   ���   ������������������������������������������������������               ���������������������               ������                  ���               ���������                           ������            ������               ���������            ���������                  ���               ���������������������������������            ���            ���            ���������������������������������               ������������������������������         ������������������������������������������������������������������������������������������������������������������������������������������      ���������������������      ������������������         ���������������������������������������������������������������������������������������������������������������   ���   ������������������������������������������������������               ������������������               ������������                                 ���������                           ������                              ������������            ������������                                 ���������������������������������                        ������            ������������������������������������            ������������������������������         ������������������������������������������������������������������������������������������������������������������������������������������         ���������������         ������������������         ���������������������������������������������������������������������������������������������������������������   ���                           ���������������������������������            ������������������               ���������������                              ���������            ������         ������������                  ������������������            ������������������                           ���������������������������������                        ������            ���������������������������������               ������������������������������         ������������������������������������������������������������������������������������������������������������������������������������������         ���������������         ������������������         ���������������������������������������������������������������������������������������                           ���������������������������   ������������������������������������            ������������               ������������������������������������            ���������������������������������������������������������������������������������������������������������������������������������            ���������������������������������                     ���������            ������������      ���������������               ������������������������������         ������������������������������������������������������������������������������������������������������������������������������������������            ������������         ���������������            ���������������������������������������������������������������������������������������   ���������������������������������������������������   ������������������������������������                                    ���������������������������������������            ���������������������������������������������������������������������������������������������������������������������������������            ���������������������������������                     ���������            ������������                                 ���������������������������������         ������������������������������������������������������������������������������������������������������������������������������������������            ������������         ���������������         ������������������������������������������������������������������������������������������   ���������������������������������������������������   ������������������������������������������                           ������������������������������������������            ������������������������������������������������������������������������������������            ���������������������������������            ���������������������������������                  ������������            ������������                              ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������         ������������         ������������            ������������������������������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������                     ���������������������������������������������            ������������������������������������������������������������������������������������            ���������������������������������            ���������������������������������               ���������������            ���������������������               ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������         ���������         ���������            ���������������������������������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������������������������������������������������������������������            ������������������������������������������������������������������������������������            ���������������������������������            ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������            ���         ���               ������������������������������������������������������������������������������������������������   ���������������������������                           ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������         ���         ������         ���������������������������������������������������������������������������������������������������                           ���   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������         ������   ���������������������������������������������������������������������������������������������������������������������������������   ���   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ������������������������������������������������������������������������������������������������������������������������������������������   ���   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             ���������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���������������������         ���         ������         ������   ������         ���         ������         ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ������������������������   ���������   ���������   ���   ������   ���������   ������������   ������   ���   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ������������������������   ������������   ������   ���   ���������   ������   ������         ������   ���   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���������������������      ������         ���   ������   ���������   ���      ������   ���������   ������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ������������������������������������������������������������������   ������������������������������������������������������������������������������������������            ���            ���         ���������            ���   ���         ������������������������������������������������������������                        ���            ���������         ���   ���            ������������������������������������������������������������   ������   ���            ���   ���������   ���         ���������         ���   ���         ���������������������������������������������         ���      ���   ���   ���               ������   ���                  ���      ���������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������������������������   ������   ���������      ���   ���   ���������������      ������      ���   ������������������������������������������������������������   ������   ���������   ���   ������   ���������������   ���������   ������   ������������������������������������������������������������   ������   ���   ������   ���   ���         ������   ���������������      ���������   ���      ������������������������������������������   ���������   ������   ���   ���               ������   ���                  ���   ������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������         ������            ���������������������������������������������������������������������������������   ������   ���         ������         ������������      ���������      ���   ������������������������������������������������������������   ������   ���      ������            ������������      ���������   ������   ������������������������������������������������������������            ���   ������   ���         ���   ������   ������������������   ���������   ���      ������������������������������������������         ���      ���         ���   ���   ���                     ���                  ���������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������   ������   ���   ������������������������������������������������������������������������������������������   ������   ���            ���   ���   ���������   ���      ���������   ���   ������������������������������������������������������������   ������   ���   ���   ���            ���������         ���������         ���������������������������������������������������������������   ������   ���            ���      ������   ������   ������������         ���������         ���������������������������������������������         ���   ������   ���������������������������������������������������������   ������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������   ������   ���   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������   ���      ���      ���   ���������������������������������������������������������������                                                                                                                     ���������������������                                                                                                                  ���������������������������                                                                                                                              ���                                                                                                                                       ���������������������������   ���������������������������������������������������   ���������������������������������������������������      ���������������   ������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ���������������������������   ������������������������������������������������������������������������������������������������������������������������   ���   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������   ���������������������������������������������������   ������������������������������������������������������������                  ���������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ���������������������������   ������������������������������������������������������������������������������������������������������������������������   ���   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������   ���������������������������������������������������   ���������������������������������������������������         ������������������      ���������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ���������������������������   ������������������������������������������������������������������������������������������������������������������������   ���   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������   ���������������������������������������������������   ���������������������������������������������      ���������������������������������      ���������������������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ���������������������������   ������������������������������������������������������������������������������������������������������������������������   ���   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������   ���������������������������������������������������   ���������������������������������������      ���������������������������������������������   ������������������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ���������������������������   ������������������������������������������������������������������������������������������������������������������������   ���   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������   ���������������������������������������������������   ������������������������������������   ������������������������������������������������������   ���������������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ���������������������������   ������������������������������������������������������������������������������������������������������������������������   ���   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������   ���������������������������������������������������   ������������������������������������   ���������������������������������������������������������   ������������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ���������������������������   ������������������������������������������������������������������������������������������������������������������������   ���   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������   ���������������������������������������������������   ���������������������������������   ������������������������������������������������������������   ������������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ���������������������������   ������������������������������������������������������������������������������������������������������������������������   ���   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������   ���������������������������������������������������   ������������������������������   ������������������������������������������������������������������   ���������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ���������������������������   ������������������������������������������������������������������������������������������������������������������������   ���   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������   ���������������������������������������������������   ������������������������������   ������������������������������������������������������������������   ���������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ���������������������������   ������������������������������������������������������������������������������������������������������������������������   ���   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������   ���������������������������                           ������������������������������   ������������������������������������������������������������������   ���������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ���������������������������   ������������������������������������������������������������������������������������������������������������������������   ���   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������                           ���   ���������������������������������������������������   ������������������������������������������������������������������������   ������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ���������������������������   ������������������������������������������������������������������������������������������������������������������������   ���   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���   ���������������������������������������������������   ������������������������������������������������������������������������   ������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ���������������������������   ������������������������������������������������������������������������������������������������������������������������   ���   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���   ���������������������������������������������������   ������������������������������������������������������������������������   ������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ���������������������������   ������������������������������������������������������������������������������������������������������������������������   ���   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���   ������������������������������������������������������   ������������������������������������������������������������������   ���������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ���������������������������   ������������������������������������������������������������������������������������������������������������������������   ���   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���   ������������������������������������������������������   ������������������������������������������������������������������   ���������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ���������������������������                                                                                                                              ���   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���   ������������������������������������������������������   ���������������������������������������������������������������   ������������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���                           ���������������������������������   ������������������������������������������������������������   ������������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������                           ���������������������������   ������������������������������������   ������������������������������������������������������   ���������������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������   ���������������������������������������������������   ������������������������������������   ������������������������������������������������������   ���������������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������   ���������������������������������������������������   ���������������������������������������   ������������������������������������������������   ������������������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������   ���������������������������������������������������   ������������������������������������������         ������������������������������         ���������������������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������   ���������������������������������������������������   ���������������������������������������������������         ������������         ������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������   ���������������������������������������������������   ������������������������������������������������������������            ���������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������   ���������������������������                           ���������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������                           ���   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���                           ���������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������                           ���������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������   ���������������������������   ���������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                       ���������������������������   ���������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������   ���������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������������������������������������������������������������������������������������������   ���������������������   ������������������������������������������������������������������������������������������������������������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���������������������������                           ���������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                     ���������������������                                                                                                                  ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                           ���   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������------BUILD07.30
----             CDL3 ���D;  ����PVBM`����  ������������h$1��1$h